** sch_path: /foss/designs/Transmission-Gate/xschem/transmission_gate.sch
**.subckt transmission_gate VDD OUT IN CONT VSS CONT_N
*.opin OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.ipin CONT
*.ipin CONT_N
XM2 IN CONT OUT VSS sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=M m=M
XM11 IN CONT_N OUT VDD sky130_fd_pr__pfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=M m=M
**.ends
.end
